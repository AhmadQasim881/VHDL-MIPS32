------------------------------------------------------------------------
-- File:           Instruction_Memory.vhdl
-- author: 	    implementing microprocessor in FBGA team
-- Description:    This is an implementation of a Instruction_Memory 
--                 behavioral architecture.
------------------------------------------------------------------------

--Library'
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.std_logic_unsigned.all;
use IEEE.NUMERIC_STD.ALL;

--Entity

entity Instruction_Memory is
port (
 ReadAddress: in std_logic_vector(31 downto 0);
 instruction: out  std_logic_vector(31 downto 0)
);
end Instruction_Memory;



--Architecture
architecture Behavioral of Instruction_Memory is


signal rom_addr: std_logic_vector(7 downto 0);
 type ROM_type is array (0 to 255 ) of std_logic_vector(31 downto 0);
 constant rom_data: ROM_type:=(

"11001100000010000000000000000000",  --LoadI @t0,@zero,0
"11001100000010010000000000000000",  --LoadI @t1,@zero,0
"11001100000100000000000000001010",  --LoadI @s0,@zero,10
"11001100000100010000000100001101",  --LoadI @s1,@zero,269
"00010010001000000000000000001011",  --beq @s1,@zero,L2
"00000010001100000101000000000110",  --Div @t2,@s1,@s0
"00000001010100000101100000101000",  --Mul @t3,@t2,@s0
"00000010001010110100100000100010",  --Sub @t1,@s1,@t3
"00000001000010010100000000100000",  --Add @t0,@t0,@t1
"00000010001100001000100000000110",  --Div @s1,@s1,@s0
"00001000000000000000000000000100",  --Jump L1
"00000001000000001011100000100000",  --Add @s7,@t0,@zero
"00000000000000000000000000000000",   --Noth
"00000000000000000000000000000000",   --Noth
"00000000000000000000000000000000",   --Noth
"00000000000000000000000000000000",   --Noth
"00000000000000000000000000000000",   --Noth
"00000000000000000000000000000000",   --Noth
"00000000000000000000000000000000",   --Noth
"00000000000000000000000000000000",   --Noth
"00000000000000000000000000000000",   --Noth
"00000000000000000000000000000000",   --Noth
"00000000000000000000000000000000",   --Noth
"00000000000000000000000000000000",   --Noth
"00000000000000000000000000000000",   --Noth
"00000000000000000000000000000000",   --Noth
"00000000000000000000000000000000",   --Noth
"00000000000000000000000000000000",   --Noth
"00000000000000000000000000000000",   --Noth
"00000000000000000000000000000000",   --Noth
"00000000000000000000000000000000",   --Noth
"00000000000000000000000000000000",   --Noth
"00000000000000000000000000000000",   --Noth
"00000000000000000000000000000000",   --Noth
"00000000000000000000000000000000",   --Noth
"00000000000000000000000000000000",   --Noth
"00000000000000000000000000000000",   --Noth
"00000000000000000000000000000000",   --Noth
"00000000000000000000000000000000",   --Noth
"00000000000000000000000000000000",   --Noth
"00000000000000000000000000000000",   --Noth
"00000000000000000000000000000000",   --Noth
"00000000000000000000000000000000",   --Noth
"00000000000000000000000000000000",   --Noth
"00000000000000000000000000000000",   --Noth
"00000000000000000000000000000000",   --Noth
"00000000000000000000000000000000",   --Noth
"00000000000000000000000000000000",   --Noth
"00000000000000000000000000000000",   --Noth
"00000000000000000000000000000000",   --Noth
"00000000000000000000000000000000",   --Noth
"00000000000000000000000000000000",   --Noth
"00000000000000000000000000000000",   --Noth
"00000000000000000000000000000000",   --Noth
"00000000000000000000000000000000",   --Noth
"00000000000000000000000000000000",   --Noth
"00000000000000000000000000000000",   --Noth
"00000000000000000000000000000000",   --Noth
"00000000000000000000000000000000",   --Noth
"00000000000000000000000000000000",   --Noth
"00000000000000000000000000000000",   --Noth
"00000000000000000000000000000000",   --Noth
"00000000000000000000000000000000",   --Noth
"00000000000000000000000000000000",   --Noth
"00000000000000000000000000000000",   --Noth
"00000000000000000000000000000000",   --Noth
"00000000000000000000000000000000",   --Noth
"00000000000000000000000000000000",   --Noth
"00000000000000000000000000000000",   --Noth
"00000000000000000000000000000000",   --Noth
"00000000000000000000000000000000",   --Noth
"00000000000000000000000000000000",   --Noth
"00000000000000000000000000000000",   --Noth
"00000000000000000000000000000000",   --Noth
"00000000000000000000000000000000",   --Noth
"00000000000000000000000000000000",   --Noth
"00000000000000000000000000000000",   --Noth
"00000000000000000000000000000000",   --Noth
"00000000000000000000000000000000",   --Noth
"00000000000000000000000000000000",   --Noth
"00000000000000000000000000000000",   --Noth
"00000000000000000000000000000000",   --Noth
"00000000000000000000000000000000",   --Noth
"00000000000000000000000000000000",   --Noth
"00000000000000000000000000000000",   --Noth
"00000000000000000000000000000000",   --Noth
"00000000000000000000000000000000",   --Noth
"00000000000000000000000000000000",   --Noth
"00000000000000000000000000000000",   --Noth
"00000000000000000000000000000000",   --Noth
"00000000000000000000000000000000",   --Noth
"00000000000000000000000000000000",   --Noth
"00000000000000000000000000000000",   --Noth
"00000000000000000000000000000000",   --Noth
"00000000000000000000000000000000",   --Noth
"00000000000000000000000000000000",   --Noth
"00000000000000000000000000000000",   --Noth
"00000000000000000000000000000000",   --Noth
"00000000000000000000000000000000",   --Noth
"00000000000000000000000000000000",   --Noth
"00000000000000000000000000000000",   --Noth
"00000000000000000000000000000000",   --Noth
"00000000000000000000000000000000",   --Noth
"00000000000000000000000000000000",   --Noth
"00000000000000000000000000000000",   --Noth
"00000000000000000000000000000000",   --Noth
"00000000000000000000000000000000",   --Noth
"00000000000000000000000000000000",   --Noth
"00000000000000000000000000000000",   --Noth
"00000000000000000000000000000000",   --Noth
"00000000000000000000000000000000",   --Noth
"00000000000000000000000000000000",   --Noth
"00000000000000000000000000000000",   --Noth
"00000000000000000000000000000000",   --Noth
"00000000000000000000000000000000",   --Noth
"00000000000000000000000000000000",   --Noth
"00000000000000000000000000000000",   --Noth
"00000000000000000000000000000000",   --Noth
"00000000000000000000000000000000",   --Noth
"00000000000000000000000000000000",   --Noth
"00000000000000000000000000000000",   --Noth
"00000000000000000000000000000000",   --Noth
"00000000000000000000000000000000",   --Noth
"00000000000000000000000000000000",   --Noth
"00000000000000000000000000000000",   --Noth
"00000000000000000000000000000000",   --Noth
"00000000000000000000000000000000",   --Noth
"00000000000000000000000000000000",   --Noth
"00000000000000000000000000000000",   --Noth
"00000000000000000000000000000000",   --Noth
"00000000000000000000000000000000",   --Noth
"00000000000000000000000000000000",   --Noth
"00000000000000000000000000000000",   --Noth
"00000000000000000000000000000000",   --Noth
"00000000000000000000000000000000",   --Noth
"00000000000000000000000000000000",   --Noth
"00000000000000000000000000000000",   --Noth
"00000000000000000000000000000000",   --Noth
"00000000000000000000000000000000",   --Noth
"00000000000000000000000000000000",   --Noth
"00000000000000000000000000000000",   --Noth
"00000000000000000000000000000000",   --Noth
"00000000000000000000000000000000",   --Noth
"00000000000000000000000000000000",   --Noth
"00000000000000000000000000000000",   --Noth
"00000000000000000000000000000000",   --Noth
"00000000000000000000000000000000",   --Noth
"00000000000000000000000000000000",   --Noth
"00000000000000000000000000000000",   --Noth
"00000000000000000000000000000000",   --Noth
"00000000000000000000000000000000",   --Noth
"00000000000000000000000000000000",   --Noth
"00000000000000000000000000000000",   --Noth
"00000000000000000000000000000000",   --Noth
"00000000000000000000000000000000",   --Noth
"00000000000000000000000000000000",   --Noth
"00000000000000000000000000000000",   --Noth
"00000000000000000000000000000000",   --Noth
"00000000000000000000000000000000",   --Noth
"00000000000000000000000000000000",   --Noth
"00000000000000000000000000000000",   --Noth
"00000000000000000000000000000000",   --Noth
"00000000000000000000000000000000",   --Noth
"00000000000000000000000000000000",   --Noth
"00000000000000000000000000000000",   --Noth
"00000000000000000000000000000000",   --Noth
"00000000000000000000000000000000",   --Noth
"00000000000000000000000000000000",   --Noth
"00000000000000000000000000000000",   --Noth
"00000000000000000000000000000000",   --Noth
"00000000000000000000000000000000",   --Noth
"00000000000000000000000000000000",   --Noth
"00000000000000000000000000000000",   --Noth
"00000000000000000000000000000000",   --Noth
"00000000000000000000000000000000",   --Noth
"00000000000000000000000000000000",   --Noth
"00000000000000000000000000000000",   --Noth
"00000000000000000000000000000000",   --Noth
"00000000000000000000000000000000",   --Noth
"00000000000000000000000000000000",   --Noth
"00000000000000000000000000000000",   --Noth
"00000000000000000000000000000000",   --Noth
"00000000000000000000000000000000",   --Noth
"00000000000000000000000000000000",   --Noth
"00000000000000000000000000000000",   --Noth
"00000000000000000000000000000000",   --Noth
"00000000000000000000000000000000",   --Noth
"00000000000000000000000000000000",   --Noth
"00000000000000000000000000000000",   --Noth
"00000000000000000000000000000000",   --Noth
"00000000000000000000000000000000",   --Noth
"00000000000000000000000000000000",   --Noth
"00000000000000000000000000000000",   --Noth
"00000000000000000000000000000000",   --Noth
"00000000000000000000000000000000",   --Noth
"00000000000000000000000000000000",   --Noth
"00000000000000000000000000000000",   --Noth
"00000000000000000000000000000000",   --Noth
"00000000000000000000000000000000",   --Noth
"00000000000000000000000000000000",   --Noth
"00000000000000000000000000000000",   --Noth
"00000000000000000000000000000000",   --Noth
"00000000000000000000000000000000",   --Noth
"00000000000000000000000000000000",   --Noth
"00000000000000000000000000000000",   --Noth
"00000000000000000000000000000000",   --Noth
"00000000000000000000000000000000",   --Noth
"00000000000000000000000000000000",   --Noth
"00000000000000000000000000000000",   --Noth
"00000000000000000000000000000000",   --Noth
"00000000000000000000000000000000",   --Noth
"00000000000000000000000000000000",   --Noth
"00000000000000000000000000000000",   --Noth
"00000000000000000000000000000000",   --Noth
"00000000000000000000000000000000",   --Noth
"00000000000000000000000000000000",   --Noth
"00000000000000000000000000000000",   --Noth
"00000000000000000000000000000000",   --Noth
"00000000000000000000000000000000",   --Noth
"00000000000000000000000000000000",   --Noth
"00000000000000000000000000000000",   --Noth
"00000000000000000000000000000000",   --Noth
"00000000000000000000000000000000",   --Noth
"00000000000000000000000000000000",   --Noth
"00000000000000000000000000000000",   --Noth
"00000000000000000000000000000000",   --Noth
"00000000000000000000000000000000",   --Noth
"00000000000000000000000000000000",   --Noth
"00000000000000000000000000000000",   --Noth
"00000000000000000000000000000000",   --Noth
"00000000000000000000000000000000",   --Noth
"00000000000000000000000000000000",   --Noth
"00000000000000000000000000000000",   --Noth
"00000000000000000000000000000000",   --Noth
"00000000000000000000000000000000",   --Noth
"00000000000000000000000000000000",   --Noth
"00000000000000000000000000000000",   --Noth
"00000000000000000000000000000000",   --Noth
"00000000000000000000000000000000",   --Noth
"00000000000000000000000000000000",   --Noth
"00000000000000000000000000000000",   --Noth
"00000000000000000000000000000000",   --Noth
"00000000000000000000000000000000",   --Noth
"00000000000000000000000000000000",   --Noth
"00000000000000000000000000000000",   --Noth
"00000000000000000000000000000000",   --Noth
"00000000000000000000000000000000",   --Noth
"00000000000000000000000000000000",   --Noth
"00000000000000000000000000000000",   --Noth
"00000000000000000000000000000000",   --Noth
"00000000000000000000000000000000",   --Noth
"00000000000000000000000000000000",   --Noth
"00000000000000000000000000000000",   --Noth
"00000000000000000000000000000000",   --Noth
"00000000000000000000000000000000",   --Noth
"00000000000000000000000000000000"    --Noth
);
begin
  
  rom_addr<=ReadAddress(9 downto 2);
  instruction <= rom_data(to_integer(unsigned(rom_addr))) when (to_integer(unsigned(ReadAddress))<1024) else x"00000000";

end Behavioral;
