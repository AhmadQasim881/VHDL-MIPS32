------------------------------------------------------------------------
-- File:           Instruction_Memory.vhdl
-- author: 	    implementing microprocessor in FBGA team
-- Description:    This is an implementation of a Instruction_Memory 
--                 behavioral architecture.
------------------------------------------------------------------------

--Library'
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.std_logic_unsigned.all;
use IEEE.NUMERIC_STD.ALL;

--Entity

entity Instruction_Memory is
port (
 ReadAddress: in std_logic_vector(31 downto 0);
 instruction: out  std_logic_vector(31 downto 0)
);
end Instruction_Memory;



--Architecture
architecture Behavioral of Instruction_Memory is


signal rom_addr: std_logic_vector(7 downto 0);
 type ROM_type is array (0 to 255 ) of std_logic_vector(31 downto 0);
 constant rom_data: ROM_type:=(

"11001100000111010000000000000000",  --LoadI @sp,@zero,0
"00001000000000000000000000110100",  --Jump main
"11001111101111010000000000000001",  --Push
"11001100000010000000000000000000",  --LoadI @t0,@zero,0
"10101111101010001111111111111111",  --Store @t0,@sp,-1
"11001100100100100000000000000000",  --LoadI @s2,@a0,0
"11001100000100110000000000000000",  --LoadI @s3,@zero,0
"01010010011100100000000001001010",  --blt @s3,@s2,Lable0
"10001111101000101111111111111111",  --Load @v0,@sp,-1
"11010011101111010000000000000001",  --Pop
"11001011111000000000000000000000",  --Jr @ra
"11010011101111010000000000000001",  --Pop
"11001011111000000000000000000000",  --Jr @ra
"10101111101111110000000000000000",  --Store @ra,@sp,0
"11001111101111010000000000000001",  --Push
"10101111101001000000000000000000",  --Store @a0,@sp,0
"11001111101111010000000000000001",  --Push
"11001100100001000000000000000000",  --LoadI @a0,@a0,0
"10001000000000000000000000000010",  --Jal reverseDigits
"11010011101111010000000000000001",  --Pop
"10001111101001000000000000000000",  --Load @a0,@sp,0
"11010011101111010000000000000001",  --Pop
"10001111101111110000000000000000",  --Load @ra,@sp,0
"11001100010001000000000000000000",  --LoadI @a0,@v0,0
"10101111101111110000000000000000",  --Store @ra,@sp,0
"11001111101111010000000000000001",  --Push
"10101111101001000000000000000000",  --Store @a0,@sp,0
"11001111101111010000000000000001",  --Push
"11001100101001000000000000000000",  --LoadI @a0,@a1,0
"10001000000000000000000000000010",  --Jal reverseDigits
"11010011101111010000000000000001",  --Pop
"10001111101001000000000000000000",  --Load @a0,@sp,0
"11010011101111010000000000000001",  --Pop
"10001111101111110000000000000000",  --Load @ra,@sp,0
"11001100010001010000000000000000",  --LoadI @a1,@v0,0
"11001111101111010000000000000001",  --Push
"11001111101111010000000000000001",  --Push
"11001100000010000000000000000000",  --LoadI @t0,@zero,0
"10101111101010001111111111111111",  --Store @t0,@sp,-1
"11001100100010000000000000000000",  --LoadI @t0,@a0,0
"10101111101010001111111111111110",  --Store @t0,@sp,-2
"10001111101101001111111111111110",  --Load @s4,@sp,-2
"11001100101101010000000000000000",  --LoadI @s5,@a1,0
"01010010100101010000000001011000",  --blt @s4,@s5,Lable4
"00010010100101010000000001011000",  --beq @s4,@s5,Lable4
"10001111101000101111111111111111",  --Load @v0,@sp,-1
"11010011101111010000000000000001",  --Pop
"11010011101111010000000000000001",  --Pop
"11001011111000000000000000000000",  --Jr @ra
"11010011101111010000000000000001",  --Pop
"11010011101111010000000000000001",  --Pop
"11001011111000000000000000000000",  --Jr @ra
"11001111101111010000000000000001",  --Push
"10101111101111110000000000000000",  --Store @ra,@sp,0
"11001111101111010000000000000001",  --Push
"10101111101001000000000000000000",  --Store @a0,@sp,0
"11001111101111010000000000000001",  --Push
"11001100000001000000000000000000",  --LoadI @a0,@zero,0
"10101111101001010000000000000000",  --Store @a1,@sp,0
"11001111101111010000000000000001",  --Push
"11001100000001010000000000010011",  --LoadI @a1,@zero,19
"10001000000000000000000000001101",  --Jal add_from_x_to_y
"11010011101111010000000000000001",  --Pop
"10001111101001010000000000000000",  --Load @a1,@sp,0
"11010011101111010000000000000001",  --Pop
"10001111101001000000000000000000",  --Load @a0,@sp,0
"11010011101111010000000000000001",  --Pop
"10001111101111110000000000000000",  --Load @ra,@sp,0
"10101111101000101111111111111111",  --Store @v0,@sp,-1
"10001111101100001111111111111111",  --Load @s0,@sp,-1
"11001110000010000000000000000000",  --AddI @t0,@s0,0
"10101111101010001111111111111111",  --Store @t0,@sp,-1
"11010011101111010000000000000001",  --Pop
"00001000000000000000000001001001",  --Jump end-labe
"10001111101100001111111111111111",  --Load @s0,@sp,-1
"11001100000000010000000000001010",  --LoadI @at,@zero,10
"00000000001100000100000000101000",  --Mul @t0,@at,@s0
"11001100000000010000000000001010",  --LoadI @at,@zero,10
"00000000100000010100100000000110",  --Div @t1,@a0,@at
"11001100000000010000000000001010",  --LoadI @at,@zero,10
"00000000001010010100100000101000",  --Mul @t1,@at,@t1
"00000000100010010100100000100010",  --Sub @t1,@a0,@t1
"00000001000010010100000000100000",  --Add @t0,@t0,@t1
"10101111101010001111111111111111",  --Store @t0,@sp,-1
"11001100000000010000000000001010",  --LoadI @at,@zero,10
"00000000100000010100000000000110",  --Div @t0,@a0,@at
"11001101000001000000000000000000",  --LoadI @a0,@t0,0
"00001000000000000000000000000101",  --Jump Lable1
"10001111101100001111111111111111",  --Load @s0,@sp,-1
"10001111101100011111111111111110",  --Load @s1,@sp,-2
"00000010000100010100000000100000",  --Add @t0,@s0,@s1
"10101111101010001111111111111111",  --Store @t0,@sp,-1
"10001111101100001111111111111110",  --Load @s0,@sp,-2
"11001110000010000000000000000001",  --AddI @t0,@s0,1
"10101111101010001111111111111110",  --Store @t0,@sp,-2
"00001000000000000000000000101001",  --Jump Lable5
"00000000000000000000000000000000",   --Noth
"00000000000000000000000000000000",   --Noth
"00000000000000000000000000000000",   --Noth
"00000000000000000000000000000000",   --Noth
"00000000000000000000000000000000",   --Noth
"00000000000000000000000000000000",   --Noth
"00000000000000000000000000000000",   --Noth
"00000000000000000000000000000000",   --Noth
"00000000000000000000000000000000",   --Noth
"00000000000000000000000000000000",   --Noth
"00000000000000000000000000000000",   --Noth
"00000000000000000000000000000000",   --Noth
"00000000000000000000000000000000",   --Noth
"00000000000000000000000000000000",   --Noth
"00000000000000000000000000000000",   --Noth
"00000000000000000000000000000000",   --Noth
"00000000000000000000000000000000",   --Noth
"00000000000000000000000000000000",   --Noth
"00000000000000000000000000000000",   --Noth
"00000000000000000000000000000000",   --Noth
"00000000000000000000000000000000",   --Noth
"00000000000000000000000000000000",   --Noth
"00000000000000000000000000000000",   --Noth
"00000000000000000000000000000000",   --Noth
"00000000000000000000000000000000",   --Noth
"00000000000000000000000000000000",   --Noth
"00000000000000000000000000000000",   --Noth
"00000000000000000000000000000000",   --Noth
"00000000000000000000000000000000",   --Noth
"00000000000000000000000000000000",   --Noth
"00000000000000000000000000000000",   --Noth
"00000000000000000000000000000000",   --Noth
"00000000000000000000000000000000",   --Noth
"00000000000000000000000000000000",   --Noth
"00000000000000000000000000000000",   --Noth
"00000000000000000000000000000000",   --Noth
"00000000000000000000000000000000",   --Noth
"00000000000000000000000000000000",   --Noth
"00000000000000000000000000000000",   --Noth
"00000000000000000000000000000000",   --Noth
"00000000000000000000000000000000",   --Noth
"00000000000000000000000000000000",   --Noth
"00000000000000000000000000000000",   --Noth
"00000000000000000000000000000000",   --Noth
"00000000000000000000000000000000",   --Noth
"00000000000000000000000000000000",   --Noth
"00000000000000000000000000000000",   --Noth
"00000000000000000000000000000000",   --Noth
"00000000000000000000000000000000",   --Noth
"00000000000000000000000000000000",   --Noth
"00000000000000000000000000000000",   --Noth
"00000000000000000000000000000000",   --Noth
"00000000000000000000000000000000",   --Noth
"00000000000000000000000000000000",   --Noth
"00000000000000000000000000000000",   --Noth
"00000000000000000000000000000000",   --Noth
"00000000000000000000000000000000",   --Noth
"00000000000000000000000000000000",   --Noth
"00000000000000000000000000000000",   --Noth
"00000000000000000000000000000000",   --Noth
"00000000000000000000000000000000",   --Noth
"00000000000000000000000000000000",   --Noth
"00000000000000000000000000000000",   --Noth
"00000000000000000000000000000000",   --Noth
"00000000000000000000000000000000",   --Noth
"00000000000000000000000000000000",   --Noth
"00000000000000000000000000000000",   --Noth
"00000000000000000000000000000000",   --Noth
"00000000000000000000000000000000",   --Noth
"00000000000000000000000000000000",   --Noth
"00000000000000000000000000000000",   --Noth
"00000000000000000000000000000000",   --Noth
"00000000000000000000000000000000",   --Noth
"00000000000000000000000000000000",   --Noth
"00000000000000000000000000000000",   --Noth
"00000000000000000000000000000000",   --Noth
"00000000000000000000000000000000",   --Noth
"00000000000000000000000000000000",   --Noth
"00000000000000000000000000000000",   --Noth
"00000000000000000000000000000000",   --Noth
"00000000000000000000000000000000",   --Noth
"00000000000000000000000000000000",   --Noth
"00000000000000000000000000000000",   --Noth
"00000000000000000000000000000000",   --Noth
"00000000000000000000000000000000",   --Noth
"00000000000000000000000000000000",   --Noth
"00000000000000000000000000000000",   --Noth
"00000000000000000000000000000000",   --Noth
"00000000000000000000000000000000",   --Noth
"00000000000000000000000000000000",   --Noth
"00000000000000000000000000000000",   --Noth
"00000000000000000000000000000000",   --Noth
"00000000000000000000000000000000",   --Noth
"00000000000000000000000000000000",   --Noth
"00000000000000000000000000000000",   --Noth
"00000000000000000000000000000000",   --Noth
"00000000000000000000000000000000",   --Noth
"00000000000000000000000000000000",   --Noth
"00000000000000000000000000000000",   --Noth
"00000000000000000000000000000000",   --Noth
"00000000000000000000000000000000",   --Noth
"00000000000000000000000000000000",   --Noth
"00000000000000000000000000000000",   --Noth
"00000000000000000000000000000000",   --Noth
"00000000000000000000000000000000",   --Noth
"00000000000000000000000000000000",   --Noth
"00000000000000000000000000000000",   --Noth
"00000000000000000000000000000000",   --Noth
"00000000000000000000000000000000",   --Noth
"00000000000000000000000000000000",   --Noth
"00000000000000000000000000000000",   --Noth
"00000000000000000000000000000000",   --Noth
"00000000000000000000000000000000",   --Noth
"00000000000000000000000000000000",   --Noth
"00000000000000000000000000000000",   --Noth
"00000000000000000000000000000000",   --Noth
"00000000000000000000000000000000",   --Noth
"00000000000000000000000000000000",   --Noth
"00000000000000000000000000000000",   --Noth
"00000000000000000000000000000000",   --Noth
"00000000000000000000000000000000",   --Noth
"00000000000000000000000000000000",   --Noth
"00000000000000000000000000000000",   --Noth
"00000000000000000000000000000000",   --Noth
"00000000000000000000000000000000",   --Noth
"00000000000000000000000000000000",   --Noth
"00000000000000000000000000000000",   --Noth
"00000000000000000000000000000000",   --Noth
"00000000000000000000000000000000",   --Noth
"00000000000000000000000000000000",   --Noth
"00000000000000000000000000000000",   --Noth
"00000000000000000000000000000000",   --Noth
"00000000000000000000000000000000",   --Noth
"00000000000000000000000000000000",   --Noth
"00000000000000000000000000000000",   --Noth
"00000000000000000000000000000000",   --Noth
"00000000000000000000000000000000",   --Noth
"00000000000000000000000000000000",   --Noth
"00000000000000000000000000000000",   --Noth
"00000000000000000000000000000000",   --Noth
"00000000000000000000000000000000",   --Noth
"00000000000000000000000000000000",   --Noth
"00000000000000000000000000000000",   --Noth
"00000000000000000000000000000000",   --Noth
"00000000000000000000000000000000",   --Noth
"00000000000000000000000000000000",   --Noth
"00000000000000000000000000000000",   --Noth
"00000000000000000000000000000000",   --Noth
"00000000000000000000000000000000",   --Noth
"00000000000000000000000000000000",   --Noth
"00000000000000000000000000000000",   --Noth
"00000000000000000000000000000000",   --Noth
"00000000000000000000000000000000",   --Noth
"00000000000000000000000000000000",   --Noth
"00000000000000000000000000000000",   --Noth
"00000000000000000000000000000000",   --Noth
"00000000000000000000000000000000",   --Noth
"00000000000000000000000000000000",   --Noth
"00000000000000000000000000000000",   --Noth
"00000000000000000000000000000000"    --Noth
);
begin
  
  rom_addr<=ReadAddress(9 downto 2);
  instruction <= rom_data(to_integer(unsigned(rom_addr))) when (to_integer(unsigned(ReadAddress))<1024) else x"00000000";

end Behavioral;
